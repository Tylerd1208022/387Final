package fmradio_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "fmradio_uvm_globals.sv"
`include "fmradio_uvm_sequence.sv"
`include "fmradio_uvm_monitor.sv"
`include "fmradio_uvm_driver.sv"
`include "fmradio_uvm_agent.sv"
`include "fmradio_uvm_scoreboard.sv"
`include "fmradio_uvm_config.sv"
`include "fmradio_uvm_env.sv"
`include "fmradio_uvm_test.sv"

endpackage
