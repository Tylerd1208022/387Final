module comparator #(
    parameter DATA_WIDTH = 32
) (
    input logic [DATA_WIDTH-1:0]     Din_L,
    input logic [DATA_WIDTH-1:0]     Din_R,
    output logic [DATA_WIDTH-1:0]    Dout,
    output logic                     isGreaterEqual
);



endmodule